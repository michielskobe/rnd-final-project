-- -------------------------------------------------------------
-- 
-- File Name: biquad.vhd
-- 
-- -------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.fixed_pkg.all;

use work.axi4_audio_pkg.all;


entity biquad is
  generic (
        g_coefficient_width : integer := 27;
        g_chip_scope : string := "False"
    );
  port( 
    -- clocking
    clk : in std_logic;

    -- axi inputs
    axi_in_fwd : in t_axi4_audio_fwd;
    axi_in_bwd : out t_axi4_audio_bwd;

    -- axi outputs
    axi_out_fwd : out t_axi4_audio_fwd;
    axi_out_bwd : in t_axi4_audio_bwd

  );
end biquad;


architecture rtl of biquad is

  -------------------------------------
  -- Memory init
  -------------------------------------
  type t_coefficient_array is array (0 to 5*2**c_ID_width) of sfixed(g_coefficient_width -1 downto 0);
  signal coefficient_array : t_coefficient_array := (others => (others => '0'));

  type t_data_array is array (0 to 4*2**c_ID_width) of signed(c_audio_width -1 downto 0);
  signal data_array : t_data_array := (others => (others => '0'));


  -------------------------------------
  -- Data Input
  -------------------------------------
  signal TData_stage_1                    : signed(23 downto 0);  -- sfix24_En23
  signal TID_stage_1                      : std_logic_vector(c_ID_width -1 downto 0);

  -------------------------------------
  -- Fetch Coefficients & Previous Data
  -------------------------------------
  signal TData_stage_2                    : signed(23 downto 0);  -- sfix24_En23
  signal TID_stage_2                      : std_logic_vector(c_ID_width -1 downto 0);

  signal Prev_Delay_X_1                   : signed(23 downto 0);  -- sfix24_En23
  signal Prev_Delay_X_2                   : signed(23 downto 0);  -- sfix24_En23
  signal Prev_Delay_Y_1                   : signed(23 downto 0);  -- sfix24_En23
  signal Prev_Delay_Y_2                   : signed(23 downto 0);  -- sfix24_En23

  signal TID_b0                           : sfixed(g_coefficient_width -1 downto 0);
  signal TID_b1                           : sfixed(g_coefficient_width -1 downto 0);
  signal TID_b2                           : sfixed(g_coefficient_width -1 downto 0);
  signal TID_a1                           : sfixed(g_coefficient_width -1 downto 0);
  signal TID_a2                           : sfixed(g_coefficient_width -1 downto 0);

  
  -------------------------------------
  -- Filter
  -------------------------------------
  -- Data
  signal TData_stage_3                    : signed(23 downto 0);  -- sfix24_En23
  signal TData_stage_4                    : signed(23 downto 0);  -- sfix24_En23
  signal TID_stage_3                      : std_logic_vector(c_ID_width -1 downto 0);
  signal TID_stage_3_prev                 : std_logic_vector(c_ID_width -1 downto 0);

  signal Prev_Delay_X_1_2                 : signed(23 downto 0);  -- sfix24_En23
  signal Prev_Delay_X_2_2                 : signed(23 downto 0);  -- sfix24_En23
  signal Prev_Delay_Y_1_2                 : signed(23 downto 0);  -- sfix24_En23
  signal Prev_Delay_Y_2_2                 : signed(23 downto 0);  -- sfix24_En23

  signal Delay_X_1                        : signed(23 downto 0);  -- sfix24_En23
  signal Delay_X_2                        : signed(23 downto 0);  -- sfix24_En23
  signal Delay_Y_1                        : signed(23 downto 0);  -- sfix24_En23
  signal Delay_Y_2                        : signed(23 downto 0);  -- sfix24_En23

  signal Delay_X_1_muxed                  : signed(23 downto 0);  -- sfix24_En23
  signal Delay_X_2_muxed                  : signed(23 downto 0);  -- sfix24_En23
  signal Delay_Y_1_muxed                  : signed(23 downto 0);  -- sfix24_En23
  signal Delay_Y_2_muxed                  : signed(23 downto 0);  -- sfix24_En23

  -- Coefficients
  signal b0_signed                        : signed(26 downto 0);  -- sfix27_En23
  signal b1_signed                        : signed(26 downto 0);  -- sfix27_En23
  signal b2_signed                        : signed(26 downto 0);  -- sfix27_En23
  signal a1_signed                        : signed(26 downto 0);  -- sfix27_En23
  signal a2_signed                        : signed(26 downto 0);  -- sfix27_En23

  signal Product1_mul_temp                : signed(50 downto 0);  -- sfix51_En46
  signal Product1_out1                    : signed(26 downto 0);  -- sfix27_En23
  signal Product2_mul_temp                : signed(50 downto 0);  -- sfix51_En46
  signal Product2_out1                    : signed(26 downto 0);  -- sfix27_En23
  signal Product3_mul_temp                : signed(50 downto 0);  -- sfix51_En46
  signal Product3_out1                    : signed(26 downto 0);  -- sfix27_En23
  signal Product4_mul_temp                : signed(50 downto 0);  -- sfix51_En46
  signal Product4_out1                    : signed(26 downto 0);  -- sfix27_En23
  signal Data_Type_Conversion_out1        : signed(23 downto 0);  -- sfix24_En23
  signal Product5_mul_temp                : signed(50 downto 0);  -- sfix51_En46
  signal Product5_out1                    : signed(26 downto 0);  -- sfix27_En23
  signal Sum2_add_cast                    : signed(31 downto 0);  -- sfix32_En23
  signal Sum2_add_cast_1                  : signed(31 downto 0);  -- sfix32_En23
  signal Sum2_out1                        : signed(31 downto 0);  -- sfix32_En23
  signal Sum1_stage2_add_cast             : signed(31 downto 0);  -- sfix32_En23
  signal Sum1_stage2_add_temp             : signed(31 downto 0);  -- sfix32_En23
  signal Sum1_op_stage1                   : signed(32 downto 0);  -- sfix33_En23
  signal Sum1_stage3_add_cast             : signed(31 downto 0);  -- sfix32_En23
  signal Sum1_stage3_add_cast_1           : signed(31 downto 0);  -- sfix32_En23
  signal Sum1_out1                        : signed(31 downto 0);  -- sfix32_En23
  signal Sum4_add_cast                    : signed(31 downto 0);  -- sfix32_En23
  signal Sum4_out1                        : signed(31 downto 0);  -- sfix32_En23


  -------------------------------------
  -- Control flow
  -------------------------------------
  signal pipe_startup : integer range 0 to 4 := 4;

   
BEGIN

  -------------------------------------
  -- Data Input
  -------------------------------------
  data_input_process : process (clk)
  begin
    if rising_edge(clk) then
      if axi_in_fwd.TValid = '1' and axi_out_bwd.TReady = '1' then
        TData_stage_1 <= signed(axi_in_fwd.TData);
        TID_stage_1 <= axi_in_fwd.TID;
      end if;
    end if;
  end process data_input_process;


  -------------------------------------
  -- Fetch Coefficients & Previous Data
  -------------------------------------
  fetch_process : process (clk)
  begin
    if rising_edge(clk) then
      if axi_in_fwd.TValid = '1' and axi_out_bwd.TReady = '1' then

        TData_stage_2 <= TData_stage_1;
        TID_stage_2 <= TID_stage_1;

        TID_b0 <= coefficient_array(5*to_integer(unsigned(TID_stage_1)));
        TID_b1 <= coefficient_array(5*to_integer(unsigned(TID_stage_1))+1);
        TID_b2 <= coefficient_array(5*to_integer(unsigned(TID_stage_1))+2);
        TID_a1 <= coefficient_array(5*to_integer(unsigned(TID_stage_1))+3);
        TID_a2 <= coefficient_array(5*to_integer(unsigned(TID_stage_1))+4);

        Prev_Delay_X_1 <= data_array(4*to_integer(unsigned(TID_stage_1)));
        Prev_Delay_X_2 <= data_array(4*to_integer(unsigned(TID_stage_1))+1);
        Prev_Delay_Y_1 <= data_array(4*to_integer(unsigned(TID_stage_1))+2);
        Prev_Delay_Y_2 <= data_array(4*to_integer(unsigned(TID_stage_1))+3);

      end if;
    end if;
  end process fetch_process;

  -------------------------------------
  -- Filter
  -------------------------------------
  filter_process : process (clk)
  begin
    if rising_edge(clk) then
      if axi_in_fwd.TValid = '1' and axi_out_bwd.TReady = '1' then

        -- Input Data
        TData_stage_3 <= TData_stage_2;
        TID_stage_3 <= TID_stage_2;
        TID_stage_3_prev <= TID_stage_3;

        Prev_Delay_X_1_2 <= Prev_Delay_X_1;
        Prev_Delay_X_2_2 <= Prev_Delay_X_2;
        Prev_Delay_Y_1_2 <= Prev_Delay_Y_1;
        Prev_Delay_Y_2_2 <= Prev_Delay_Y_2;

        -- Z^-1
        Delay_X_1 <= TData_stage_3;
        Delay_X_2 <= Delay_X_1_muxed;
        Delay_Y_1 <= Data_Type_Conversion_out1;
        Delay_Y_2 <= Delay_Y_1_muxed;

        -- Move Coefficients to Filter
        b0_signed <= signed(TID_b0);
        b1_signed <= signed(TID_b1);
        b2_signed <= signed(TID_b2);
        a1_signed <= signed(TID_a1);
        a2_signed <= signed(TID_a2);

        -- Move Data from Filter
        data_array(4*to_integer(unsigned(TID_stage_3_prev)))   <= Delay_X_1;
        data_array(4*to_integer(unsigned(TID_stage_3_prev))+1) <= Delay_X_2;
        data_array(4*to_integer(unsigned(TID_stage_3_prev))+2) <= Delay_Y_1;
        data_array(4*to_integer(unsigned(TID_stage_3_prev))+3) <= Delay_Y_2;

      end if;
    end if;
  end process filter_process;


  mux : process (all)
  begin

    -- Mux to choose between the current Delay if TID = TID_prev or the Prev_Delay if TID != TID_prev
    if TID_stage_3 /= TID_stage_3_prev then
      Delay_X_1_muxed <= Prev_Delay_X_1_2;
      Delay_X_2_muxed <= Prev_Delay_X_2_2;
      Delay_Y_1_muxed <= Prev_Delay_Y_1_2;
      Delay_Y_2_muxed <= Prev_Delay_Y_2_2;
    else
      Delay_X_1_muxed <= Delay_X_1;
      Delay_X_2_muxed <= Delay_X_2;
      Delay_Y_1_muxed <= Delay_Y_1;
      Delay_Y_2_muxed <= Delay_Y_2;
    end if;
    
  end process mux;
  

  -- Product 1
  Product1_mul_temp <= TData_stage_3 * b0_signed;
  Product1_out1 <= Product1_mul_temp(49 downto 23);
  
  -- Product 2
  Product2_mul_temp <= Delay_X_1_muxed * b1_signed;
  Product2_out1 <= Product2_mul_temp(49 downto 23);

  -- Product 3
  Product3_mul_temp <= Delay_X_2_muxed * b2_signed;
  Product3_out1 <= Product3_mul_temp(49 downto 23);

  -- Product 4
  Product4_mul_temp <= Delay_Y_1_muxed * a1_signed;
  Product4_out1 <= Product4_mul_temp(49 downto 23);

  -- Product 5
  Product5_mul_temp <= Delay_Y_2_muxed * a2_signed;
  Product5_out1 <= Product5_mul_temp(49 downto 23);

  -- Sum of Product 3 & Product 5
  Sum2_add_cast <= resize(Product3_out1, 32);
  Sum2_add_cast_1 <= resize(Product5_out1, 32);
  Sum2_out1 <= Sum2_add_cast + Sum2_add_cast_1;

  -- Sum of Product 2 & Product 4 & Sum 2
  Sum1_stage2_add_cast <= resize(Product2_out1, 32);
  Sum1_stage2_add_temp <= Sum1_stage2_add_cast + Sum2_out1;
  Sum1_op_stage1 <= resize(Sum1_stage2_add_temp, 33);
  Sum1_stage3_add_cast <= Sum1_op_stage1(31 downto 0);
  Sum1_stage3_add_cast_1 <= resize(Product4_out1, 32);
  Sum1_out1 <= Sum1_stage3_add_cast + Sum1_stage3_add_cast_1;

  -- Sum of Product 1 & Sum 1
  Sum4_add_cast <= resize(Product1_out1, 32);
  Sum4_out1 <= Sum4_add_cast + Sum1_out1;

  -- Output conversion
  Data_Type_Conversion_out1 <= Sum4_out1(23 downto 0);
  TData_stage_4 <= Data_Type_Conversion_out1;

  -------------------------------------
  -- Output Data
  -------------------------------------
  data_output_process : process (clk)
  begin
    if rising_edge(clk) then
      if axi_in_fwd.TValid = '1' and axi_out_bwd.TReady = '1' then

        axi_out_fwd.TData <= std_logic_vector(TData_stage_4);
        axi_out_fwd.TID   <= TID_stage_3;

      end if;
    end if;
  end process data_output_process;


  -------------------------------------
  -- Control flow
  -------------------------------------
  -- we are ready if the module behind us is ready
  axi_in_bwd.TReady <= axi_out_bwd.TReady;

  p_ctrl_flow : process (clk)
  begin
      if rising_edge(clk) then
          if axi_in_fwd.TValid = '1' and axi_out_bwd.TReady = '1' then

              if pipe_startup = 0 then
                pipe_startup <= pipe_startup;
              else
                pipe_startup <= pipe_startup - 1;
              end if;

          end if;
      end if;
  end process;


  p_valid : process (all)
  begin

      if pipe_startup = 0 then
          axi_out_fwd.TValid <= axi_in_fwd.TValid;
      else
          axi_out_fwd.TValid <= '0';
      end if;

  end process;


END rtl;
